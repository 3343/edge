////
// @file This file is part of EDGE.
//
// @author Alexander Breuer (anbreuer AT ucsd.edu)
//
// @section LICENSE
// Copyright (c) 2017, Regents of the University of California
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without modification, are permitted provided that the following conditions are met:
//
// 1. Redistributions of source code must retain the above copyright notice, this list of conditions and the following disclaimer.
//
// 2. Redistributions in binary form must reproduce the above copyright notice, this list of conditions and the following disclaimer in the documentation and/or other materials provided with the distribution.
//
// 3. Neither the name of the copyright holder nor the names of its contributors may be used to endorse or promote products derived from this software without specific prior written permission.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// @section DESCRIPTION
// netCDF-template for benchmarks using kinematic sources
////
netcdf {
types:
  compound Vector3 {
    double x;
    double y;
    double z;
  };

  compound Subfault_units {
    string tinit;
    string timestep;
    string mu;
    string area;
    string tan1;
    string tan2;
    string normal;
  };

  compound Subfault {
    double tinit;
    double timestep;
    double mu;
    double area;
    Vector3 tan1;
    Vector3 tan2;
    Vector3 normal;
  };

dimensions:
        source = TEMPLATE_N_SRC;

variables:
        Vector3 centres(source);
                centres:units = "m";
        Subfault subfaults(source) ;
                Subfault_units subfaults:units = {"s", "s", "pascal", "m^2", "m", "m", "m"};
data:
  centres   = TEMPLATE_CENTERS;
  subfaults = TEMPLATE_SUBFAULTS;
}
